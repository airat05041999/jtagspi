//////////////////////////////////////////////////
//~:(
//@module: Spi_interface_test.sv
//@author: Yafizov Airat
//@date: 15.12.2021
//@version: 1.0.0
//@description: testbench 
//~:)
//////////////////////////////////////////////////
`timescale 10 ns/10 ns
//////////////////////////////////////////////////
module spi_top_test;

//////////////////////////////////////////////////
//Local signals
//////////////////////////////////////////////////

logic clk;
logic rst;
logic miso;

//////////////////////////////////////////////////
//Tested module
//////////////////////////////////////////////////

spi_top spi_top_inst (
    .clk(clk), .rst(rst),
    .miso(miso)
    );

//////////////////////////////////////////////////
//Test
//////////////////////////////////////////////////

initial
    begin
        rst = 1;
        #10;
        rst = 0;
    end

//////////////////////////////////////////////////
//clk
//////////////////////////////////////////////////

initial                                                
    begin                                                  
        clk=0;
        forever #5 clk=~clk;
    end

initial                                                
    begin                                                  
        miso=1;
        forever #10 miso=~miso;
    end

endmodule
